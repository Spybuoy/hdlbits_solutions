module top_module (
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);//

    wire c_wire, c;
    add16 inst1(a[15:0], b[15:0], 1'b0, sum[15:0], c_wire);
    add16 inst2(a[31:16], b[31:16], c_wire, sum[31:16], c);

    
endmodule

module add1 ( input a, input b, input cin,   output sum, output cout );

// Full adder module here
    assign {cout, sum} = a+b+cin;

endmodule
