module fa(input a,input b,input cin,output sum,output cout);
    assign {cout, sum} = a+b+cin;
endmodule
    

module top_module( 
    input [99:0] a, b,
    input cin,
    output [99:0] cout,
    output [99:0] sum );
	
    generate
    	genvar i;
        for(i=0;i<100;i=i+1)
            begin:loop
                if(i==0)
                    begin
                        fa inst1(.a(a[i]), .b(b[i]), .cin(cin),.sum(sum[i]), .cout(cout[i]));
                    end
                else
                    begin
                        fa inst2(.a(a[i]), .b(b[i]), .cin(cout[i-1]),.sum(sum[i]), .cout(cout[i]));
                    end
            end
    endgenerate
endmodule
